library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity toplevel is
end toplevel;

architecture Behavioral of toplevel is

begin


end Behavioral;

